// soc1.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc1 (
		inout  wire        accelerometer_spi_I2C_SDAT,      // accelerometer_spi.I2C_SDAT
		output wire        accelerometer_spi_I2C_SCLK,      //                  .I2C_SCLK
		output wire        accelerometer_spi_G_SENSOR_CS_N, //                  .G_SENSOR_CS_N
		input  wire        accelerometer_spi_G_SENSOR_INT,  //                  .G_SENSOR_INT
		input  wire        clk_clk,                         //               clk.clk
		output wire [3:0]  hex0_export,                     //              hex0.export
		output wire [3:0]  hex1_export,                     //              hex1.export
		output wire [3:0]  hex2_export,                     //              hex2.export
		output wire [3:0]  hex3_export,                     //              hex3.export
		output wire [3:0]  hex4_export,                     //              hex4.export
		output wire [3:0]  hex5_export,                     //              hex5.export
		input  wire [1:0]  key_export,                      //               key.export
		output wire [9:0]  ledr_export,                     //              ledr.export
		input  wire        reset_reset_n,                   //             reset.reset_n
		output wire        sdram_clk_clk,                   //         sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                 //        sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                   //                  .ba
		output wire        sdram_wire_cas_n,                //                  .cas_n
		output wire        sdram_wire_cke,                  //                  .cke
		output wire        sdram_wire_cs_n,                 //                  .cs_n
		inout  wire [15:0] sdram_wire_dq,                   //                  .dq
		output wire [1:0]  sdram_wire_dqm,                  //                  .dqm
		output wire        sdram_wire_ras_n,                //                  .ras_n
		output wire        sdram_wire_we_n,                 //                  .we_n
		input  wire [9:0]  sw_export,                       //                sw.export
		output wire        vga_out_CLK,                     //           vga_out.CLK
		output wire        vga_out_HS,                      //                  .HS
		output wire        vga_out_VS,                      //                  .VS
		output wire        vga_out_BLANK,                   //                  .BLANK
		output wire        vga_out_SYNC,                    //                  .SYNC
		output wire [3:0]  vga_out_R,                       //                  .R
		output wire [3:0]  vga_out_G,                       //                  .G
		output wire [3:0]  vga_out_B                        //                  .B
	);

	wire         video_change_alpha_0_avalon_apply_alpha_source_valid;                                  // video_change_alpha_0:stream_out_valid -> video_alpha_blender_0:foreground_valid
	wire  [39:0] video_change_alpha_0_avalon_apply_alpha_source_data;                                   // video_change_alpha_0:stream_out_data -> video_alpha_blender_0:foreground_data
	wire         video_change_alpha_0_avalon_apply_alpha_source_ready;                                  // video_alpha_blender_0:foreground_ready -> video_change_alpha_0:stream_out_ready
	wire         video_change_alpha_0_avalon_apply_alpha_source_startofpacket;                          // video_change_alpha_0:stream_out_startofpacket -> video_alpha_blender_0:foreground_startofpacket
	wire         video_change_alpha_0_avalon_apply_alpha_source_endofpacket;                            // video_change_alpha_0:stream_out_endofpacket -> video_alpha_blender_0:foreground_endofpacket
	wire         video_alpha_blender_0_avalon_blended_source_valid;                                     // video_alpha_blender_0:output_valid -> video_dual_clock_buffer_0:stream_in_valid
	wire  [29:0] video_alpha_blender_0_avalon_blended_source_data;                                      // video_alpha_blender_0:output_data -> video_dual_clock_buffer_0:stream_in_data
	wire         video_alpha_blender_0_avalon_blended_source_ready;                                     // video_dual_clock_buffer_0:stream_in_ready -> video_alpha_blender_0:output_ready
	wire         video_alpha_blender_0_avalon_blended_source_startofpacket;                             // video_alpha_blender_0:output_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	wire         video_alpha_blender_0_avalon_blended_source_endofpacket;                               // video_alpha_blender_0:output_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	wire         charbuff_avalon_char_source_valid;                                                     // charbuff:stream_valid -> video_change_alpha_0:stream_in_valid
	wire  [39:0] charbuff_avalon_char_source_data;                                                      // charbuff:stream_data -> video_change_alpha_0:stream_in_data
	wire         charbuff_avalon_char_source_ready;                                                     // video_change_alpha_0:stream_in_ready -> charbuff:stream_ready
	wire         charbuff_avalon_char_source_startofpacket;                                             // charbuff:stream_startofpacket -> video_change_alpha_0:stream_in_startofpacket
	wire         charbuff_avalon_char_source_endofpacket;                                               // charbuff:stream_endofpacket -> video_change_alpha_0:stream_in_endofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;                               // video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	wire  [29:0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;                                // video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;                               // video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;                       // video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;                         // video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire         pixelbuff_avalon_pixel_source_valid;                                                   // pixelbuff:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire   [7:0] pixelbuff_avalon_pixel_source_data;                                                    // pixelbuff:stream_data -> video_rgb_resampler_0:stream_in_data
	wire         pixelbuff_avalon_pixel_source_ready;                                                   // video_rgb_resampler_0:stream_in_ready -> pixelbuff:stream_ready
	wire         pixelbuff_avalon_pixel_source_startofpacket;                                           // pixelbuff:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         pixelbuff_avalon_pixel_source_endofpacket;                                             // pixelbuff:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;                                         // video_rgb_resampler_0:stream_out_valid -> video_scaler_0:stream_in_valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                                          // video_rgb_resampler_0:stream_out_data -> video_scaler_0:stream_in_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;                                         // video_scaler_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;                                 // video_rgb_resampler_0:stream_out_startofpacket -> video_scaler_0:stream_in_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;                                   // video_rgb_resampler_0:stream_out_endofpacket -> video_scaler_0:stream_in_endofpacket
	wire         pll_c0_clk;                                                                            // pll:c0 -> [accelerometer_spi_0:clk, avalon_st_adapter:in_clk_0_clk, charbuff:clk, cpu:clk, hex0:clk, hex1:clk, hex2:clk, hex3:clk, hex4:clk, hex5:clk, irq_mapper:clk, jtag_uart:clk, key:clk, ledr:clk, mm_interconnect_0:pll_c0_clk, pixelbuff:clk, ram:clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, sw:clk, sysid_qsys_0:clock, timer_0:clk, video_alpha_blender_0:clk, video_change_alpha_0:clk, video_dual_clock_buffer_0:clk_stream_in, video_rgb_resampler_0:clk, video_scaler_0:clk]
	wire         pll_c2_clk;                                                                            // pll:c2 -> [rst_controller_003:clk, rst_controller_004:clk, video_dual_clock_buffer_0:clk_stream_out, video_vga_controller_0:clk]
	wire         pixelbuff_avalon_pixel_dma_master_waitrequest;                                         // mm_interconnect_0:pixelbuff_avalon_pixel_dma_master_waitrequest -> pixelbuff:master_waitrequest
	wire   [7:0] pixelbuff_avalon_pixel_dma_master_readdata;                                            // mm_interconnect_0:pixelbuff_avalon_pixel_dma_master_readdata -> pixelbuff:master_readdata
	wire  [31:0] pixelbuff_avalon_pixel_dma_master_address;                                             // pixelbuff:master_address -> mm_interconnect_0:pixelbuff_avalon_pixel_dma_master_address
	wire         pixelbuff_avalon_pixel_dma_master_read;                                                // pixelbuff:master_read -> mm_interconnect_0:pixelbuff_avalon_pixel_dma_master_read
	wire         pixelbuff_avalon_pixel_dma_master_readdatavalid;                                       // mm_interconnect_0:pixelbuff_avalon_pixel_dma_master_readdatavalid -> pixelbuff:master_readdatavalid
	wire         pixelbuff_avalon_pixel_dma_master_lock;                                                // pixelbuff:master_arbiterlock -> mm_interconnect_0:pixelbuff_avalon_pixel_dma_master_lock
	wire  [31:0] cpu_data_master_readdata;                                                              // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                                           // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                                           // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                                               // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                                            // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                                  // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                                         // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                                                 // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                             // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                                       // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                                    // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                                                        // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                                           // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                                  // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_ram_s1_chipselect;                                                   // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                                                     // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire  [14:0] mm_interconnect_0_ram_s1_address;                                                      // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                                                   // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;                                                        // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                                                    // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                                                        // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire   [7:0] mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata;    // accelerometer_spi_0:readdata -> mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata
	wire         mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest; // accelerometer_spi_0:waitrequest -> mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest
	wire   [0:0] mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address;     // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address -> accelerometer_spi_0:address
	wire         mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read;        // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read -> accelerometer_spi_0:read
	wire   [0:0] mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable;  // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable -> accelerometer_spi_0:byteenable
	wire         mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write;       // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write -> accelerometer_spi_0:write
	wire   [7:0] mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata;   // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata -> accelerometer_spi_0:writedata
	wire         mm_interconnect_0_charbuff_avalon_char_buffer_slave_chipselect;                        // mm_interconnect_0:charbuff_avalon_char_buffer_slave_chipselect -> charbuff:buf_chipselect
	wire   [7:0] mm_interconnect_0_charbuff_avalon_char_buffer_slave_readdata;                          // charbuff:buf_readdata -> mm_interconnect_0:charbuff_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_charbuff_avalon_char_buffer_slave_waitrequest;                       // charbuff:buf_waitrequest -> mm_interconnect_0:charbuff_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_charbuff_avalon_char_buffer_slave_address;                           // mm_interconnect_0:charbuff_avalon_char_buffer_slave_address -> charbuff:buf_address
	wire         mm_interconnect_0_charbuff_avalon_char_buffer_slave_read;                              // mm_interconnect_0:charbuff_avalon_char_buffer_slave_read -> charbuff:buf_read
	wire   [0:0] mm_interconnect_0_charbuff_avalon_char_buffer_slave_byteenable;                        // mm_interconnect_0:charbuff_avalon_char_buffer_slave_byteenable -> charbuff:buf_byteenable
	wire         mm_interconnect_0_charbuff_avalon_char_buffer_slave_write;                             // mm_interconnect_0:charbuff_avalon_char_buffer_slave_write -> charbuff:buf_write
	wire   [7:0] mm_interconnect_0_charbuff_avalon_char_buffer_slave_writedata;                         // mm_interconnect_0:charbuff_avalon_char_buffer_slave_writedata -> charbuff:buf_writedata
	wire         mm_interconnect_0_charbuff_avalon_char_control_slave_chipselect;                       // mm_interconnect_0:charbuff_avalon_char_control_slave_chipselect -> charbuff:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_charbuff_avalon_char_control_slave_readdata;                         // charbuff:ctrl_readdata -> mm_interconnect_0:charbuff_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_charbuff_avalon_char_control_slave_address;                          // mm_interconnect_0:charbuff_avalon_char_control_slave_address -> charbuff:ctrl_address
	wire         mm_interconnect_0_charbuff_avalon_char_control_slave_read;                             // mm_interconnect_0:charbuff_avalon_char_control_slave_read -> charbuff:ctrl_read
	wire   [3:0] mm_interconnect_0_charbuff_avalon_char_control_slave_byteenable;                       // mm_interconnect_0:charbuff_avalon_char_control_slave_byteenable -> charbuff:ctrl_byteenable
	wire         mm_interconnect_0_charbuff_avalon_char_control_slave_write;                            // mm_interconnect_0:charbuff_avalon_char_control_slave_write -> charbuff:ctrl_write
	wire  [31:0] mm_interconnect_0_charbuff_avalon_char_control_slave_writedata;                        // mm_interconnect_0:charbuff_avalon_char_control_slave_writedata -> charbuff:ctrl_writedata
	wire  [31:0] mm_interconnect_0_pixelbuff_avalon_control_slave_readdata;                             // pixelbuff:slave_readdata -> mm_interconnect_0:pixelbuff_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pixelbuff_avalon_control_slave_address;                              // mm_interconnect_0:pixelbuff_avalon_control_slave_address -> pixelbuff:slave_address
	wire         mm_interconnect_0_pixelbuff_avalon_control_slave_read;                                 // mm_interconnect_0:pixelbuff_avalon_control_slave_read -> pixelbuff:slave_read
	wire   [3:0] mm_interconnect_0_pixelbuff_avalon_control_slave_byteenable;                           // mm_interconnect_0:pixelbuff_avalon_control_slave_byteenable -> pixelbuff:slave_byteenable
	wire         mm_interconnect_0_pixelbuff_avalon_control_slave_write;                                // mm_interconnect_0:pixelbuff_avalon_control_slave_write -> pixelbuff:slave_write
	wire  [31:0] mm_interconnect_0_pixelbuff_avalon_control_slave_writedata;                            // mm_interconnect_0:pixelbuff_avalon_control_slave_writedata -> pixelbuff:slave_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                                // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                             // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata;                     // video_rgb_resampler_0:slave_readdata -> mm_interconnect_0:video_rgb_resampler_0_avalon_rgb_slave_readdata
	wire         mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read;                         // mm_interconnect_0:video_rgb_resampler_0_avalon_rgb_slave_read -> video_rgb_resampler_0:slave_read
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                                 // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                                  // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                                        // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                                     // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                                     // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                                         // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                                            // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                                      // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                                           // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                                       // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                                              // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                                               // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                                                  // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                                                 // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                                             // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                                 // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                                   // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                                // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                                    // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                       // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                                 // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                              // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                      // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                                  // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_0_s1_chipselect;                                               // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                                 // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                                  // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                                    // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                                                // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_hex0_s1_chipselect;                                                  // mm_interconnect_0:hex0_s1_chipselect -> hex0:chipselect
	wire  [31:0] mm_interconnect_0_hex0_s1_readdata;                                                    // hex0:readdata -> mm_interconnect_0:hex0_s1_readdata
	wire   [2:0] mm_interconnect_0_hex0_s1_address;                                                     // mm_interconnect_0:hex0_s1_address -> hex0:address
	wire         mm_interconnect_0_hex0_s1_write;                                                       // mm_interconnect_0:hex0_s1_write -> hex0:write_n
	wire  [31:0] mm_interconnect_0_hex0_s1_writedata;                                                   // mm_interconnect_0:hex0_s1_writedata -> hex0:writedata
	wire         mm_interconnect_0_hex1_s1_chipselect;                                                  // mm_interconnect_0:hex1_s1_chipselect -> hex1:chipselect
	wire  [31:0] mm_interconnect_0_hex1_s1_readdata;                                                    // hex1:readdata -> mm_interconnect_0:hex1_s1_readdata
	wire   [2:0] mm_interconnect_0_hex1_s1_address;                                                     // mm_interconnect_0:hex1_s1_address -> hex1:address
	wire         mm_interconnect_0_hex1_s1_write;                                                       // mm_interconnect_0:hex1_s1_write -> hex1:write_n
	wire  [31:0] mm_interconnect_0_hex1_s1_writedata;                                                   // mm_interconnect_0:hex1_s1_writedata -> hex1:writedata
	wire         mm_interconnect_0_hex2_s1_chipselect;                                                  // mm_interconnect_0:hex2_s1_chipselect -> hex2:chipselect
	wire  [31:0] mm_interconnect_0_hex2_s1_readdata;                                                    // hex2:readdata -> mm_interconnect_0:hex2_s1_readdata
	wire   [2:0] mm_interconnect_0_hex2_s1_address;                                                     // mm_interconnect_0:hex2_s1_address -> hex2:address
	wire         mm_interconnect_0_hex2_s1_write;                                                       // mm_interconnect_0:hex2_s1_write -> hex2:write_n
	wire  [31:0] mm_interconnect_0_hex2_s1_writedata;                                                   // mm_interconnect_0:hex2_s1_writedata -> hex2:writedata
	wire         mm_interconnect_0_hex3_s1_chipselect;                                                  // mm_interconnect_0:hex3_s1_chipselect -> hex3:chipselect
	wire  [31:0] mm_interconnect_0_hex3_s1_readdata;                                                    // hex3:readdata -> mm_interconnect_0:hex3_s1_readdata
	wire   [2:0] mm_interconnect_0_hex3_s1_address;                                                     // mm_interconnect_0:hex3_s1_address -> hex3:address
	wire         mm_interconnect_0_hex3_s1_write;                                                       // mm_interconnect_0:hex3_s1_write -> hex3:write_n
	wire  [31:0] mm_interconnect_0_hex3_s1_writedata;                                                   // mm_interconnect_0:hex3_s1_writedata -> hex3:writedata
	wire         mm_interconnect_0_hex4_s1_chipselect;                                                  // mm_interconnect_0:hex4_s1_chipselect -> hex4:chipselect
	wire  [31:0] mm_interconnect_0_hex4_s1_readdata;                                                    // hex4:readdata -> mm_interconnect_0:hex4_s1_readdata
	wire   [2:0] mm_interconnect_0_hex4_s1_address;                                                     // mm_interconnect_0:hex4_s1_address -> hex4:address
	wire         mm_interconnect_0_hex4_s1_write;                                                       // mm_interconnect_0:hex4_s1_write -> hex4:write_n
	wire  [31:0] mm_interconnect_0_hex4_s1_writedata;                                                   // mm_interconnect_0:hex4_s1_writedata -> hex4:writedata
	wire         mm_interconnect_0_hex5_s1_chipselect;                                                  // mm_interconnect_0:hex5_s1_chipselect -> hex5:chipselect
	wire  [31:0] mm_interconnect_0_hex5_s1_readdata;                                                    // hex5:readdata -> mm_interconnect_0:hex5_s1_readdata
	wire   [2:0] mm_interconnect_0_hex5_s1_address;                                                     // mm_interconnect_0:hex5_s1_address -> hex5:address
	wire         mm_interconnect_0_hex5_s1_write;                                                       // mm_interconnect_0:hex5_s1_write -> hex5:write_n
	wire  [31:0] mm_interconnect_0_hex5_s1_writedata;                                                   // mm_interconnect_0:hex5_s1_writedata -> hex5:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                                                      // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [2:0] mm_interconnect_0_sw_s1_address;                                                       // mm_interconnect_0:sw_s1_address -> sw:address
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                                                     // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [2:0] mm_interconnect_0_key_s1_address;                                                      // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_ledr_s1_chipselect;                                                  // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                                                    // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [2:0] mm_interconnect_0_ledr_s1_address;                                                     // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_write;                                                       // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                                                   // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire         irq_mapper_receiver0_irq;                                                              // accelerometer_spi_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                              // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                              // timer_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                                                           // irq_mapper:sender_irq -> cpu:irq
	wire         video_scaler_0_avalon_scaler_source_valid;                                             // video_scaler_0:stream_out_valid -> avalon_st_adapter:in_0_valid
	wire  [29:0] video_scaler_0_avalon_scaler_source_data;                                              // video_scaler_0:stream_out_data -> avalon_st_adapter:in_0_data
	wire         video_scaler_0_avalon_scaler_source_ready;                                             // avalon_st_adapter:in_0_ready -> video_scaler_0:stream_out_ready
	wire   [3:0] video_scaler_0_avalon_scaler_source_channel;                                           // video_scaler_0:stream_out_channel -> avalon_st_adapter:in_0_channel
	wire         video_scaler_0_avalon_scaler_source_startofpacket;                                     // video_scaler_0:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         video_scaler_0_avalon_scaler_source_endofpacket;                                       // video_scaler_0:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                                         // avalon_st_adapter:out_0_valid -> video_alpha_blender_0:background_valid
	wire  [29:0] avalon_st_adapter_out_0_data;                                                          // avalon_st_adapter:out_0_data -> video_alpha_blender_0:background_data
	wire         avalon_st_adapter_out_0_ready;                                                         // video_alpha_blender_0:background_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                                                 // avalon_st_adapter:out_0_startofpacket -> video_alpha_blender_0:background_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                                                   // avalon_st_adapter:out_0_endofpacket -> video_alpha_blender_0:background_endofpacket
	wire         rst_controller_reset_out_reset;                                                        // rst_controller:reset_out -> [accelerometer_spi_0:reset, avalon_st_adapter:in_rst_0_reset, charbuff:reset, cpu:reset_n, hex0:reset_n, hex1:reset_n, hex2:reset_n, hex3:reset_n, hex4:reset_n, hex5:reset_n, irq_mapper:reset, key:reset_n, ledr:reset_n, mm_interconnect_0:pixelbuff_reset_reset_bridge_in_reset_reset, pixelbuff:reset, ram:reset, rst_translator:in_reset, sdram:reset_n, sw:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, video_change_alpha_0:reset, video_rgb_resampler_0:reset, video_scaler_0:reset]
	wire         rst_controller_reset_out_reset_req;                                                    // rst_controller:reset_req -> [cpu:reset_req, ram:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                                    // rst_controller_001:reset_out -> [jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, video_alpha_blender_0:reset, video_dual_clock_buffer_0:reset_stream_in]
	wire         cpu_debug_reset_request_reset;                                                         // cpu:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_002_reset_out_reset;                                                    // rst_controller_002:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]
	wire         rst_controller_003_reset_out_reset;                                                    // rst_controller_003:reset_out -> video_dual_clock_buffer_0:reset_stream_out
	wire         rst_controller_004_reset_out_reset;                                                    // rst_controller_004:reset_out -> video_vga_controller_0:reset

	soc1_accelerometer_spi_0 accelerometer_spi_0 (
		.clk           (pll_c0_clk),                                                                            //                                 clk.clk
		.reset         (rst_controller_reset_out_reset),                                                        //                               reset.reset
		.address       (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address),     // avalon_accelerometer_spi_mode_slave.address
		.byteenable    (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable),  //                                    .byteenable
		.read          (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read),        //                                    .read
		.write         (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write),       //                                    .write
		.writedata     (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata),   //                                    .writedata
		.readdata      (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata),    //                                    .readdata
		.waitrequest   (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest), //                                    .waitrequest
		.irq           (irq_mapper_receiver0_irq),                                                              //                           interrupt.irq
		.I2C_SDAT      (accelerometer_spi_I2C_SDAT),                                                            //                  external_interface.export
		.I2C_SCLK      (accelerometer_spi_I2C_SCLK),                                                            //                                    .export
		.G_SENSOR_CS_N (accelerometer_spi_G_SENSOR_CS_N),                                                       //                                    .export
		.G_SENSOR_INT  (accelerometer_spi_G_SENSOR_INT)                                                         //                                    .export
	);

	soc1_charbuff charbuff (
		.clk                  (pll_c0_clk),                                                      //                       clk.clk
		.reset                (rst_controller_reset_out_reset),                                  //                     reset.reset
		.ctrl_address         (mm_interconnect_0_charbuff_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_charbuff_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_charbuff_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_charbuff_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_charbuff_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_charbuff_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_charbuff_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_charbuff_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_charbuff_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_charbuff_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_charbuff_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_charbuff_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_charbuff_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_charbuff_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_charbuff_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (charbuff_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (charbuff_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (charbuff_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (charbuff_avalon_char_source_valid),                               //                          .valid
		.stream_data          (charbuff_avalon_char_source_data)                                 //                          .data
	);

	soc1_cpu cpu (
		.clk                                 (pll_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	soc1_hex0 hex0 (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex0_export)                           // external_connection.export
	);

	soc1_hex0 hex1 (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex1_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                           // external_connection.export
	);

	soc1_hex0 hex2 (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex2_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                           // external_connection.export
	);

	soc1_hex0 hex3 (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_s1_readdata),   //                    .readdata
		.out_port   (hex3_export)                           // external_connection.export
	);

	soc1_hex0 hex4 (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex4_export)                           // external_connection.export
	);

	soc1_hex0 hex5 (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_s1_readdata),   //                    .readdata
		.out_port   (hex5_export)                           // external_connection.export
	);

	soc1_jtag_uart jtag_uart (
		.clk            (pll_c0_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	soc1_key key (
		.clk      (pll_c0_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata), //                    .readdata
		.in_port  (key_export)                         // external_connection.export
	);

	soc1_ledr ledr (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	soc1_pixelbuff pixelbuff (
		.clk                  (pll_c0_clk),                                                  //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                              //                   reset.reset
		.master_readdatavalid (pixelbuff_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixelbuff_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixelbuff_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixelbuff_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixelbuff_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixelbuff_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixelbuff_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixelbuff_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixelbuff_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixelbuff_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixelbuff_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixelbuff_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixelbuff_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixelbuff_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixelbuff_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixelbuff_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixelbuff_avalon_pixel_source_data)                           //                        .data
	);

	soc1_pll pll (
		.clk                (clk_clk),                                   //       inclk_interface.clk
		.reset              (rst_controller_002_reset_out_reset),        // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0                 (pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                             //                    c1.clk
		.c2                 (pll_c2_clk),                                //                    c2.clk
		.scandone           (),                                          //           (terminated)
		.scandataout        (),                                          //           (terminated)
		.c3                 (),                                          //           (terminated)
		.c4                 (),                                          //           (terminated)
		.areset             (1'b0),                                      //           (terminated)
		.locked             (),                                          //           (terminated)
		.phasedone          (),                                          //           (terminated)
		.phasecounterselect (3'b000),                                    //           (terminated)
		.phaseupdown        (1'b0),                                      //           (terminated)
		.phasestep          (1'b0),                                      //           (terminated)
		.scanclk            (1'b0),                                      //           (terminated)
		.scanclkena         (1'b0),                                      //           (terminated)
		.scandata           (1'b0),                                      //           (terminated)
		.configupdate       (1'b0)                                       //           (terminated)
	);

	soc1_ram ram (
		.clk        (pll_c0_clk),                          //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	soc1_sdram sdram (
		.clk            (pll_c0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	soc1_sw sw (
		.clk      (pll_c0_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_export)                         // external_connection.export
	);

	soc1_sysid_qsys_0 sysid_qsys_0 (
		.clock    (pll_c0_clk),                                            //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	soc1_timer_0 timer_0 (
		.clk        (pll_c0_clk),                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	soc1_video_alpha_blender_0 video_alpha_blender_0 (
		.clk                      (pll_c0_clk),                                                   //                    clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                           //                  reset.reset
		.foreground_data          (video_change_alpha_0_avalon_apply_alpha_source_data),          // avalon_foreground_sink.data
		.foreground_startofpacket (video_change_alpha_0_avalon_apply_alpha_source_startofpacket), //                       .startofpacket
		.foreground_endofpacket   (video_change_alpha_0_avalon_apply_alpha_source_endofpacket),   //                       .endofpacket
		.foreground_valid         (video_change_alpha_0_avalon_apply_alpha_source_valid),         //                       .valid
		.foreground_ready         (video_change_alpha_0_avalon_apply_alpha_source_ready),         //                       .ready
		.background_data          (avalon_st_adapter_out_0_data),                                 // avalon_background_sink.data
		.background_startofpacket (avalon_st_adapter_out_0_startofpacket),                        //                       .startofpacket
		.background_endofpacket   (avalon_st_adapter_out_0_endofpacket),                          //                       .endofpacket
		.background_valid         (avalon_st_adapter_out_0_valid),                                //                       .valid
		.background_ready         (avalon_st_adapter_out_0_ready),                                //                       .ready
		.output_ready             (video_alpha_blender_0_avalon_blended_source_ready),            //  avalon_blended_source.ready
		.output_data              (video_alpha_blender_0_avalon_blended_source_data),             //                       .data
		.output_startofpacket     (video_alpha_blender_0_avalon_blended_source_startofpacket),    //                       .startofpacket
		.output_endofpacket       (video_alpha_blender_0_avalon_blended_source_endofpacket),      //                       .endofpacket
		.output_valid             (video_alpha_blender_0_avalon_blended_source_valid)             //                       .valid
	);

	soc1_video_change_alpha_0 video_change_alpha_0 (
		.clk                      (pll_c0_clk),                                                   //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                               //                     reset.reset
		.stream_in_startofpacket  (charbuff_avalon_char_source_startofpacket),                    //   avalon_apply_alpha_sink.startofpacket
		.stream_in_endofpacket    (charbuff_avalon_char_source_endofpacket),                      //                          .endofpacket
		.stream_in_valid          (charbuff_avalon_char_source_valid),                            //                          .valid
		.stream_in_ready          (charbuff_avalon_char_source_ready),                            //                          .ready
		.stream_in_data           (charbuff_avalon_char_source_data),                             //                          .data
		.stream_out_ready         (video_change_alpha_0_avalon_apply_alpha_source_ready),         // avalon_apply_alpha_source.ready
		.stream_out_startofpacket (video_change_alpha_0_avalon_apply_alpha_source_startofpacket), //                          .startofpacket
		.stream_out_endofpacket   (video_change_alpha_0_avalon_apply_alpha_source_endofpacket),   //                          .endofpacket
		.stream_out_valid         (video_change_alpha_0_avalon_apply_alpha_source_valid),         //                          .valid
		.stream_out_data          (video_change_alpha_0_avalon_apply_alpha_source_data)           //                          .data
	);

	soc1_video_dual_clock_buffer_0 video_dual_clock_buffer_0 (
		.clk_stream_in            (pll_c0_clk),                                                      //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_001_reset_out_reset),                              //         reset_stream_in.reset
		.clk_stream_out           (pll_c2_clk),                                                      //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_003_reset_out_reset),                              //        reset_stream_out.reset
		.stream_in_ready          (video_alpha_blender_0_avalon_blended_source_ready),               //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_alpha_blender_0_avalon_blended_source_startofpacket),       //                        .startofpacket
		.stream_in_endofpacket    (video_alpha_blender_0_avalon_blended_source_endofpacket),         //                        .endofpacket
		.stream_in_valid          (video_alpha_blender_0_avalon_blended_source_valid),               //                        .valid
		.stream_in_data           (video_alpha_blender_0_avalon_blended_source_data),                //                        .data
		.stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data)           //                        .data
	);

	soc1_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (pll_c0_clk),                                                        //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //             reset.reset
		.stream_in_startofpacket  (pixelbuff_avalon_pixel_source_startofpacket),                       //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixelbuff_avalon_pixel_source_endofpacket),                         //                  .endofpacket
		.stream_in_valid          (pixelbuff_avalon_pixel_source_valid),                               //                  .valid
		.stream_in_ready          (pixelbuff_avalon_pixel_source_ready),                               //                  .ready
		.stream_in_data           (pixelbuff_avalon_pixel_source_data),                                //                  .data
		.slave_read               (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read),     //  avalon_rgb_slave.read
		.slave_readdata           (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata), //                  .readdata
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),                     // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),             //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),               //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),                     //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)                       //                  .data
	);

	soc1_video_scaler_0 video_scaler_0 (
		.clk                      (pll_c0_clk),                                            //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                        //                reset.reset
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (video_scaler_0_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_0_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_0_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (video_scaler_0_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (video_scaler_0_avalon_scaler_source_data),              //                     .data
		.stream_out_channel       (video_scaler_0_avalon_scaler_source_channel)            //                     .channel
	);

	soc1_video_vga_controller_0 video_vga_controller_0 (
		.clk           (pll_c2_clk),                                                      //                clk.clk
		.reset         (rst_controller_004_reset_out_reset),                              //              reset.reset
		.data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_out_CLK),                                                     // external_interface.export
		.VGA_HS        (vga_out_HS),                                                      //                   .export
		.VGA_VS        (vga_out_VS),                                                      //                   .export
		.VGA_BLANK     (vga_out_BLANK),                                                   //                   .export
		.VGA_SYNC      (vga_out_SYNC),                                                    //                   .export
		.VGA_R         (vga_out_R),                                                       //                   .export
		.VGA_G         (vga_out_G),                                                       //                   .export
		.VGA_B         (vga_out_B)                                                        //                   .export
	);

	soc1_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                       (clk_clk),                                                                               //                                               clk_0_clk.clk
		.pll_c0_clk                                                          (pll_c0_clk),                                                                            //                                                  pll_c0.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset                         (rst_controller_001_reset_out_reset),                                                    //                   jtag_uart_reset_reset_bridge_in_reset.reset
		.pixelbuff_reset_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),                                                        //                   pixelbuff_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset               (rst_controller_002_reset_out_reset),                                                    //         pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                             (cpu_data_master_address),                                                               //                                         cpu_data_master.address
		.cpu_data_master_waitrequest                                         (cpu_data_master_waitrequest),                                                           //                                                        .waitrequest
		.cpu_data_master_byteenable                                          (cpu_data_master_byteenable),                                                            //                                                        .byteenable
		.cpu_data_master_read                                                (cpu_data_master_read),                                                                  //                                                        .read
		.cpu_data_master_readdata                                            (cpu_data_master_readdata),                                                              //                                                        .readdata
		.cpu_data_master_readdatavalid                                       (cpu_data_master_readdatavalid),                                                         //                                                        .readdatavalid
		.cpu_data_master_write                                               (cpu_data_master_write),                                                                 //                                                        .write
		.cpu_data_master_writedata                                           (cpu_data_master_writedata),                                                             //                                                        .writedata
		.cpu_data_master_debugaccess                                         (cpu_data_master_debugaccess),                                                           //                                                        .debugaccess
		.cpu_instruction_master_address                                      (cpu_instruction_master_address),                                                        //                                  cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                                  (cpu_instruction_master_waitrequest),                                                    //                                                        .waitrequest
		.cpu_instruction_master_read                                         (cpu_instruction_master_read),                                                           //                                                        .read
		.cpu_instruction_master_readdata                                     (cpu_instruction_master_readdata),                                                       //                                                        .readdata
		.cpu_instruction_master_readdatavalid                                (cpu_instruction_master_readdatavalid),                                                  //                                                        .readdatavalid
		.pixelbuff_avalon_pixel_dma_master_address                           (pixelbuff_avalon_pixel_dma_master_address),                                             //                       pixelbuff_avalon_pixel_dma_master.address
		.pixelbuff_avalon_pixel_dma_master_waitrequest                       (pixelbuff_avalon_pixel_dma_master_waitrequest),                                         //                                                        .waitrequest
		.pixelbuff_avalon_pixel_dma_master_read                              (pixelbuff_avalon_pixel_dma_master_read),                                                //                                                        .read
		.pixelbuff_avalon_pixel_dma_master_readdata                          (pixelbuff_avalon_pixel_dma_master_readdata),                                            //                                                        .readdata
		.pixelbuff_avalon_pixel_dma_master_readdatavalid                     (pixelbuff_avalon_pixel_dma_master_readdatavalid),                                       //                                                        .readdatavalid
		.pixelbuff_avalon_pixel_dma_master_lock                              (pixelbuff_avalon_pixel_dma_master_lock),                                                //                                                        .lock
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address     (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address),     // accelerometer_spi_0_avalon_accelerometer_spi_mode_slave.address
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write       (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write),       //                                                        .write
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read        (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read),        //                                                        .read
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata    (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata),    //                                                        .readdata
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata   (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata),   //                                                        .writedata
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable  (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable),  //                                                        .byteenable
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest), //                                                        .waitrequest
		.charbuff_avalon_char_buffer_slave_address                           (mm_interconnect_0_charbuff_avalon_char_buffer_slave_address),                           //                       charbuff_avalon_char_buffer_slave.address
		.charbuff_avalon_char_buffer_slave_write                             (mm_interconnect_0_charbuff_avalon_char_buffer_slave_write),                             //                                                        .write
		.charbuff_avalon_char_buffer_slave_read                              (mm_interconnect_0_charbuff_avalon_char_buffer_slave_read),                              //                                                        .read
		.charbuff_avalon_char_buffer_slave_readdata                          (mm_interconnect_0_charbuff_avalon_char_buffer_slave_readdata),                          //                                                        .readdata
		.charbuff_avalon_char_buffer_slave_writedata                         (mm_interconnect_0_charbuff_avalon_char_buffer_slave_writedata),                         //                                                        .writedata
		.charbuff_avalon_char_buffer_slave_byteenable                        (mm_interconnect_0_charbuff_avalon_char_buffer_slave_byteenable),                        //                                                        .byteenable
		.charbuff_avalon_char_buffer_slave_waitrequest                       (mm_interconnect_0_charbuff_avalon_char_buffer_slave_waitrequest),                       //                                                        .waitrequest
		.charbuff_avalon_char_buffer_slave_chipselect                        (mm_interconnect_0_charbuff_avalon_char_buffer_slave_chipselect),                        //                                                        .chipselect
		.charbuff_avalon_char_control_slave_address                          (mm_interconnect_0_charbuff_avalon_char_control_slave_address),                          //                      charbuff_avalon_char_control_slave.address
		.charbuff_avalon_char_control_slave_write                            (mm_interconnect_0_charbuff_avalon_char_control_slave_write),                            //                                                        .write
		.charbuff_avalon_char_control_slave_read                             (mm_interconnect_0_charbuff_avalon_char_control_slave_read),                             //                                                        .read
		.charbuff_avalon_char_control_slave_readdata                         (mm_interconnect_0_charbuff_avalon_char_control_slave_readdata),                         //                                                        .readdata
		.charbuff_avalon_char_control_slave_writedata                        (mm_interconnect_0_charbuff_avalon_char_control_slave_writedata),                        //                                                        .writedata
		.charbuff_avalon_char_control_slave_byteenable                       (mm_interconnect_0_charbuff_avalon_char_control_slave_byteenable),                       //                                                        .byteenable
		.charbuff_avalon_char_control_slave_chipselect                       (mm_interconnect_0_charbuff_avalon_char_control_slave_chipselect),                       //                                                        .chipselect
		.cpu_debug_mem_slave_address                                         (mm_interconnect_0_cpu_debug_mem_slave_address),                                         //                                     cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                           (mm_interconnect_0_cpu_debug_mem_slave_write),                                           //                                                        .write
		.cpu_debug_mem_slave_read                                            (mm_interconnect_0_cpu_debug_mem_slave_read),                                            //                                                        .read
		.cpu_debug_mem_slave_readdata                                        (mm_interconnect_0_cpu_debug_mem_slave_readdata),                                        //                                                        .readdata
		.cpu_debug_mem_slave_writedata                                       (mm_interconnect_0_cpu_debug_mem_slave_writedata),                                       //                                                        .writedata
		.cpu_debug_mem_slave_byteenable                                      (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                                      //                                                        .byteenable
		.cpu_debug_mem_slave_waitrequest                                     (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                                     //                                                        .waitrequest
		.cpu_debug_mem_slave_debugaccess                                     (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                                     //                                                        .debugaccess
		.hex0_s1_address                                                     (mm_interconnect_0_hex0_s1_address),                                                     //                                                 hex0_s1.address
		.hex0_s1_write                                                       (mm_interconnect_0_hex0_s1_write),                                                       //                                                        .write
		.hex0_s1_readdata                                                    (mm_interconnect_0_hex0_s1_readdata),                                                    //                                                        .readdata
		.hex0_s1_writedata                                                   (mm_interconnect_0_hex0_s1_writedata),                                                   //                                                        .writedata
		.hex0_s1_chipselect                                                  (mm_interconnect_0_hex0_s1_chipselect),                                                  //                                                        .chipselect
		.hex1_s1_address                                                     (mm_interconnect_0_hex1_s1_address),                                                     //                                                 hex1_s1.address
		.hex1_s1_write                                                       (mm_interconnect_0_hex1_s1_write),                                                       //                                                        .write
		.hex1_s1_readdata                                                    (mm_interconnect_0_hex1_s1_readdata),                                                    //                                                        .readdata
		.hex1_s1_writedata                                                   (mm_interconnect_0_hex1_s1_writedata),                                                   //                                                        .writedata
		.hex1_s1_chipselect                                                  (mm_interconnect_0_hex1_s1_chipselect),                                                  //                                                        .chipselect
		.hex2_s1_address                                                     (mm_interconnect_0_hex2_s1_address),                                                     //                                                 hex2_s1.address
		.hex2_s1_write                                                       (mm_interconnect_0_hex2_s1_write),                                                       //                                                        .write
		.hex2_s1_readdata                                                    (mm_interconnect_0_hex2_s1_readdata),                                                    //                                                        .readdata
		.hex2_s1_writedata                                                   (mm_interconnect_0_hex2_s1_writedata),                                                   //                                                        .writedata
		.hex2_s1_chipselect                                                  (mm_interconnect_0_hex2_s1_chipselect),                                                  //                                                        .chipselect
		.hex3_s1_address                                                     (mm_interconnect_0_hex3_s1_address),                                                     //                                                 hex3_s1.address
		.hex3_s1_write                                                       (mm_interconnect_0_hex3_s1_write),                                                       //                                                        .write
		.hex3_s1_readdata                                                    (mm_interconnect_0_hex3_s1_readdata),                                                    //                                                        .readdata
		.hex3_s1_writedata                                                   (mm_interconnect_0_hex3_s1_writedata),                                                   //                                                        .writedata
		.hex3_s1_chipselect                                                  (mm_interconnect_0_hex3_s1_chipselect),                                                  //                                                        .chipselect
		.hex4_s1_address                                                     (mm_interconnect_0_hex4_s1_address),                                                     //                                                 hex4_s1.address
		.hex4_s1_write                                                       (mm_interconnect_0_hex4_s1_write),                                                       //                                                        .write
		.hex4_s1_readdata                                                    (mm_interconnect_0_hex4_s1_readdata),                                                    //                                                        .readdata
		.hex4_s1_writedata                                                   (mm_interconnect_0_hex4_s1_writedata),                                                   //                                                        .writedata
		.hex4_s1_chipselect                                                  (mm_interconnect_0_hex4_s1_chipselect),                                                  //                                                        .chipselect
		.hex5_s1_address                                                     (mm_interconnect_0_hex5_s1_address),                                                     //                                                 hex5_s1.address
		.hex5_s1_write                                                       (mm_interconnect_0_hex5_s1_write),                                                       //                                                        .write
		.hex5_s1_readdata                                                    (mm_interconnect_0_hex5_s1_readdata),                                                    //                                                        .readdata
		.hex5_s1_writedata                                                   (mm_interconnect_0_hex5_s1_writedata),                                                   //                                                        .writedata
		.hex5_s1_chipselect                                                  (mm_interconnect_0_hex5_s1_chipselect),                                                  //                                                        .chipselect
		.jtag_uart_avalon_jtag_slave_address                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                                 //                             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                                   //                                                        .write
		.jtag_uart_avalon_jtag_slave_read                                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                                    //                                                        .read
		.jtag_uart_avalon_jtag_slave_readdata                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                                //                                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                               //                                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),                             //                                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                              //                                                        .chipselect
		.key_s1_address                                                      (mm_interconnect_0_key_s1_address),                                                      //                                                  key_s1.address
		.key_s1_readdata                                                     (mm_interconnect_0_key_s1_readdata),                                                     //                                                        .readdata
		.ledr_s1_address                                                     (mm_interconnect_0_ledr_s1_address),                                                     //                                                 ledr_s1.address
		.ledr_s1_write                                                       (mm_interconnect_0_ledr_s1_write),                                                       //                                                        .write
		.ledr_s1_readdata                                                    (mm_interconnect_0_ledr_s1_readdata),                                                    //                                                        .readdata
		.ledr_s1_writedata                                                   (mm_interconnect_0_ledr_s1_writedata),                                                   //                                                        .writedata
		.ledr_s1_chipselect                                                  (mm_interconnect_0_ledr_s1_chipselect),                                                  //                                                        .chipselect
		.pixelbuff_avalon_control_slave_address                              (mm_interconnect_0_pixelbuff_avalon_control_slave_address),                              //                          pixelbuff_avalon_control_slave.address
		.pixelbuff_avalon_control_slave_write                                (mm_interconnect_0_pixelbuff_avalon_control_slave_write),                                //                                                        .write
		.pixelbuff_avalon_control_slave_read                                 (mm_interconnect_0_pixelbuff_avalon_control_slave_read),                                 //                                                        .read
		.pixelbuff_avalon_control_slave_readdata                             (mm_interconnect_0_pixelbuff_avalon_control_slave_readdata),                             //                                                        .readdata
		.pixelbuff_avalon_control_slave_writedata                            (mm_interconnect_0_pixelbuff_avalon_control_slave_writedata),                            //                                                        .writedata
		.pixelbuff_avalon_control_slave_byteenable                           (mm_interconnect_0_pixelbuff_avalon_control_slave_byteenable),                           //                                                        .byteenable
		.pll_pll_slave_address                                               (mm_interconnect_0_pll_pll_slave_address),                                               //                                           pll_pll_slave.address
		.pll_pll_slave_write                                                 (mm_interconnect_0_pll_pll_slave_write),                                                 //                                                        .write
		.pll_pll_slave_read                                                  (mm_interconnect_0_pll_pll_slave_read),                                                  //                                                        .read
		.pll_pll_slave_readdata                                              (mm_interconnect_0_pll_pll_slave_readdata),                                              //                                                        .readdata
		.pll_pll_slave_writedata                                             (mm_interconnect_0_pll_pll_slave_writedata),                                             //                                                        .writedata
		.ram_s1_address                                                      (mm_interconnect_0_ram_s1_address),                                                      //                                                  ram_s1.address
		.ram_s1_write                                                        (mm_interconnect_0_ram_s1_write),                                                        //                                                        .write
		.ram_s1_readdata                                                     (mm_interconnect_0_ram_s1_readdata),                                                     //                                                        .readdata
		.ram_s1_writedata                                                    (mm_interconnect_0_ram_s1_writedata),                                                    //                                                        .writedata
		.ram_s1_byteenable                                                   (mm_interconnect_0_ram_s1_byteenable),                                                   //                                                        .byteenable
		.ram_s1_chipselect                                                   (mm_interconnect_0_ram_s1_chipselect),                                                   //                                                        .chipselect
		.ram_s1_clken                                                        (mm_interconnect_0_ram_s1_clken),                                                        //                                                        .clken
		.sdram_s1_address                                                    (mm_interconnect_0_sdram_s1_address),                                                    //                                                sdram_s1.address
		.sdram_s1_write                                                      (mm_interconnect_0_sdram_s1_write),                                                      //                                                        .write
		.sdram_s1_read                                                       (mm_interconnect_0_sdram_s1_read),                                                       //                                                        .read
		.sdram_s1_readdata                                                   (mm_interconnect_0_sdram_s1_readdata),                                                   //                                                        .readdata
		.sdram_s1_writedata                                                  (mm_interconnect_0_sdram_s1_writedata),                                                  //                                                        .writedata
		.sdram_s1_byteenable                                                 (mm_interconnect_0_sdram_s1_byteenable),                                                 //                                                        .byteenable
		.sdram_s1_readdatavalid                                              (mm_interconnect_0_sdram_s1_readdatavalid),                                              //                                                        .readdatavalid
		.sdram_s1_waitrequest                                                (mm_interconnect_0_sdram_s1_waitrequest),                                                //                                                        .waitrequest
		.sdram_s1_chipselect                                                 (mm_interconnect_0_sdram_s1_chipselect),                                                 //                                                        .chipselect
		.sw_s1_address                                                       (mm_interconnect_0_sw_s1_address),                                                       //                                                   sw_s1.address
		.sw_s1_readdata                                                      (mm_interconnect_0_sw_s1_readdata),                                                      //                                                        .readdata
		.sysid_qsys_0_control_slave_address                                  (mm_interconnect_0_sysid_qsys_0_control_slave_address),                                  //                              sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                 (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                                 //                                                        .readdata
		.timer_0_s1_address                                                  (mm_interconnect_0_timer_0_s1_address),                                                  //                                              timer_0_s1.address
		.timer_0_s1_write                                                    (mm_interconnect_0_timer_0_s1_write),                                                    //                                                        .write
		.timer_0_s1_readdata                                                 (mm_interconnect_0_timer_0_s1_readdata),                                                 //                                                        .readdata
		.timer_0_s1_writedata                                                (mm_interconnect_0_timer_0_s1_writedata),                                                //                                                        .writedata
		.timer_0_s1_chipselect                                               (mm_interconnect_0_timer_0_s1_chipselect),                                               //                                                        .chipselect
		.video_rgb_resampler_0_avalon_rgb_slave_read                         (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read),                         //                  video_rgb_resampler_0_avalon_rgb_slave.read
		.video_rgb_resampler_0_avalon_rgb_slave_readdata                     (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata)                      //                                                        .readdata
	);

	soc1_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	soc1_avalon_st_adapter #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (4),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (pll_c0_clk),                                        // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                    // in_rst_0.reset
		.in_0_data           (video_scaler_0_avalon_scaler_source_data),          //     in_0.data
		.in_0_valid          (video_scaler_0_avalon_scaler_source_valid),         //         .valid
		.in_0_ready          (video_scaler_0_avalon_scaler_source_ready),         //         .ready
		.in_0_startofpacket  (video_scaler_0_avalon_scaler_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (video_scaler_0_avalon_scaler_source_endofpacket),   //         .endofpacket
		.in_0_channel        (video_scaler_0_avalon_scaler_source_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                      //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                     //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                     //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),             //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (pll_c2_clk),                         //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_c2_clk),                         //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
